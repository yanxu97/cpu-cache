library verilog;
use verilog.vl_types.all;
entity load_byte_mask_sv_unit is
end load_byte_mask_sv_unit;
