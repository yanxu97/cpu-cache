library verilog;
use verilog.vl_types.all;
entity mp0_sv_unit is
end mp0_sv_unit;
