library verilog;
use verilog.vl_types.all;
entity modifier_sv_unit is
end modifier_sv_unit;
