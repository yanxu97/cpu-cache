library verilog;
use verilog.vl_types.all;
entity cmp_sv_unit is
end cmp_sv_unit;
