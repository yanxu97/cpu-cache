library verilog;
use verilog.vl_types.all;
entity mp1_sv_unit is
end mp1_sv_unit;
