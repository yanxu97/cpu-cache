library verilog;
use verilog.vl_types.all;
entity cpu_control_sv_unit is
end cpu_control_sv_unit;
