library verilog;
use verilog.vl_types.all;
entity mp1_tb is
end mp1_tb;
