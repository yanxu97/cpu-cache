library verilog;
use verilog.vl_types.all;
entity mp0_tb is
end mp0_tb;
