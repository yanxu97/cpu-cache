library verilog;
use verilog.vl_types.all;
entity rv32i_types is
end rv32i_types;
